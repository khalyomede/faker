module faker

pub fn (currency Currency) to_code() string {
    return match currency {
        .afghani { "AFN" }
        .argentina_peso { "ARS" }
        .aruba_guilder { "AWG" }
        .australia_dollar { "AUD" }
        .bahamas_dollar { "BSD" }
        .baht { "THB" }
        .balboa { "PAB" }
        .barbados_dollar { "BBD" }
        .belarus_ruble { "BYN" }
        .belize_dollar { "BZD" }
        .bermuda_dollar { "BMD" }
        .brunei_darusalam_dollar { "BND" }
        .bolivar { "VES" }
        .boliviano { "BOB" }
        .convertible_mark { "BAM" }
        .canada_dollar { "CAD" }
        .cayman_islands_dollar { "KYD" }
        .cedi { "GHS" }
        .chile_peso { "CLP" }
        .colombia_peso { "COP" }
        .cordoba { "NIO" }
        .costa_rica_colon { "CRC" }
        .cuba_peso { "CUP" }
        .denar { "MKD" }
        .denmark_krone { "DKK" }
        .dong { "VND" }
        .dominican_republic_peso { "DOP" }
        .east_caribbean_dollar { "XCD" }
        .egypt_pound { "EGP" }
        .euro { "EUR" }
        .falkland_islands_pound { "FKP" }
        .forint { "HUF" }
        .fiji_dollar { "FJD" }
        .gibraltar_pound { "GIP" }
        .guarani { "PYG" }
        .guernsey_pound { "GGP" }
        .guyana_dollar { "GYD" }
        .hong_kong_dollar { "HKD" }
        .hryvnia { "UAH" }
        .iceland_krona { "ISK" }
        .india_rupee { "INR" }
        .iran_riyal { "IRR" }
        .isle_of_man_pound { "IMP" }
        .jamaica_dollar { "JMD" }
        .jersey_pound { "JEP" }
        .koruna { "CZK" }
        .kip { "LAK" }
        .kuna { "HRK" }
        .kyrgyzstan_som { "KGS" }
        .lebanon_pound { "LBP" }
        .lek { "ALL" }
        .lempira { "HNL" }
        .leu { "RON" }
        .lev { "BGN" }
        .liberia_dollar { "LRD" }
        .lira { "TRY" }
        .azerbaijan_manat { "AZN" }
        .mauritius_rupee { "MUR" }
        .mexico_peso { "MXN" }
        .metical { "MZN" }
        .naira { "NGN" }
        .namibia_dollar { "NAD" }
        .nepal_rupee { "NPR" }
        .netherlands_antilles_guilder { "ANG" }
        .new_taiwan_dollar { "TWD" }
        .new_zealand_dollar { "NZD" }
        .north_korea_won { "KPW" }
        .norway_krone { "NOK" }
        .oman_riyal { "OMR" }
        .pakistan_rupee { "PKR" }
        .philipine_peso { "PHP" }
        .pula { "BWP" }
        .qatar_riyal { "QAR" }
        .quetzal { "GTQ" }
        .rand { "ZAR" }
        .real { "BRL" }
        .riel { "KHR" }
        .ringgit { "MYR" }
        .rupiah { "IDR" }
        .russia_ruble { "RUB" }
        .saint_helena_pound { "SHP" }
        .saudi_arabia_riyal { "SAR" }
        .serbia_dinar { "RSD" }
        .seychelles_rupee { "SCR" }
        .shekel { "ILS" }
        .shilling { "KES" }
        .singapore_dollar { "SGD" }
        .sol { "PEN" }
        .solomon_islands_dollar { "SBD" }
        .south_korea_won { "KRW" }
        .sri_lanka_rupee { "LKR" }
        .suriname_dollar { "SRD" }
        .sweden_krona { "SEK" }
        .switzerland_franc { "CHF" }
        .syria_pound { "SYP" }
        .tenge { "KZT" }
        .trinidad_and_tobago_dollar { "TTD" }
        .tughrik { "MNT" }
        .turkmenistan_manat { "TMT" }
        .tuvalu_dollar { "TVD" }
        .united_kingdom_pound { "GBP" }
        .united_states_dollar { "USD" }
        .uruguay_peso { "UYU" }
        .uzbekistan_som { "UZS" }
        .yen { "JPY" }
        .yemen_riyal { "YER" }
        .yuan { "CNY" }
        .zimbabwe_dollar { "ZWL" }
        .zloty { "PLN" }
    }
}
