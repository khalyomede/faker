module faker

pub enum Country {
    afghanistan
    albania
    algeria
    andorra
    angola
    antigua_and_barbuda
    argentina
    armenia
    australia
    austria
    azerbaijan
    bahamas
    bahrain
    bangladesh
    barbados
    belarus
    belgium
    belize
    benin
    bhutan
    bolivia
    bosnia_and_herzegovina
    botswana
    brazil
    brunei
    bulgaria
    burkina_faso
    burundi
    cabo_verde
    cambodia
    cameroon
    canada
    central_african_republic
    chad
    chile
    china
    colombia
    comoros
    congo
    costa_rica
    croatia
    cuba
    cyprus
    czech_republic
    democratic_republic_of_the_congo
    denmark
    djibouti
    dominica
    dominican_republic
    ecuador
    egypt
    el_salvador
    equatorial_guinea
    eritrea
    estonia
    eswatini
    ethiopia
    fiji
    finland
    france
    gabon
    gambia
    georgia
    germany
    ghana
    greece
    grenada
    guatemala
    guinea
    guinea_bissau
    guyana
    haiti
    holy_see
    honduras
    hungary
    iceland
    india
    indonesia
    iran
    iraq
    ireland
    israel
    italy
    ivory_coast
    jamaica
    japan
    jordan
    kazakhstan
    kenya
    kiribati
    kosovo
    kuwait
    kyrgyzstan
    laos
    latvia
    lebanon
    lesotho
    liberia
    libya
    liechtenstein
    lithuania
    luxembourg
    madagascar
    malawi
    malaysia
    maldives
    mali
    malta
    marshall_islands
    mauritania
    mauritius
    mexico
    micronesia
    moldova
    monaco
    mongolia
    montenegro
    morocco
    mozambique
    myanmar
    namibia
    nauru
    nepal
    netherlands
    new_zealand
    nicaragua
    niger
    nigeria
    north_korea
    north_macedonia
    norway
    oman
    pakistan
    palau
    palestine
    panama
    papua_new_guinea
    paraguay
    peru
    philippines
    poland
    portugal
    qatar
    romania
    russia
    rwanda
    saint_kitts_and_nevis
    saint_lucia
    saint_vincent_and_the_grenadines
    samoa
    san_marino
    sao_tome_and_principe
    saudi_arabia
    senegal
    serbia
    seychelles
    sierra_leone
    singapore
    slovakia
    slovenia
    solomon_islands
    somalia
    south_africa
    south_korea
    south_sudan
    spain
    sri_lanka
    sudan
    suriname
    sweden
    switzerland
    syria
    taiwan
    tajikistan
    tanzania
    thailand
    timor_leste
    togo
    tonga
    trinidad_and_tobago
    tunisia
    turkey
    turkmenistan
    tuvalu
    uganda
    ukraine
    united_arab_emirates
    united_kingdom
    united_states
    uruguay
    uzbekistan
    vanuatu
    venezuela
    vietnam
    yemen
    zambia
    zimbabwe
}
