module faker

pub enum Lang {
    en
}
