module faker

pub struct RandomLineInFileParameters {
    file   string
    not_tied_to_lang bool
}
