module faker

pub struct FakerU8BetweenParameters {
    pub:
        min u8
        max u8
}
