module faker

pub struct FakerI32BetweenParameters {
    pub:
        min i32
        max i32
}
