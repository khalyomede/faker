module faker

pub struct FakerU64BetweenParameters {
    pub:
        min u64
        max u64
}
