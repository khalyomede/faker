module faker

pub struct FakerF32BetweenParameters {
    pub:
        min f32
        max f32
}
