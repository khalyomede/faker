module faker

pub fn (currency Currency) to_symbol() string {
    return match currency {
        .afghani { "؋" }
        .argentina_peso { "\$" }
        .aruba_guilder { "ƒ" }
        .australia_dollar { "\$" }
        .bahamas_dollar { "\$" }
        .baht { "฿" }
        .balboa { "B/." }
        .barbados_dollar { "\$" }
        .belarus_ruble { "Br" }
        .belize_dollar { "BZ$" }
        .bermuda_dollar { "\$" }
        .brunei_darusalam_dollar { "\$" }
        .bolivar { "Bs." }
        .boliviano { "Bs" }
        .convertible_mark { "КМ" }
        .canada_dollar { "\$" }
        .cayman_islands_dollar { "\$" }
        .cedi { "₵" }
        .chile_peso { "\$" }
        .colombia_peso { "\$" }
        .cordoba { "C$" }
        .costa_rica_colon { "₡" }
        .cuba_peso { "₱" }
        .denar { "ден" }
        .denmark_krone { "kr" }
        .dong { "₫" }
        .dominican_republic_peso { "RD$" }
        .east_caribbean_dollar { "\$" }
        .egypt_pound { "£" }
        .euro { "€" }
        .falkland_islands_pound { "£" }
        .forint { "Ft" }
        .fiji_dollar { "\$" }
        .gibraltar_pound { "£" }
        .guarani { "₲" }
        .guernsey_pound { "£" }
        .guyana_dollar { "\$" }
        .hong_kong_dollar { "\$" }
        .hryvnia { "₴" }
        .iceland_krona { "kr" }
        .india_rupee { "₹" }
        .iran_riyal { "﷼" }
        .isle_of_man_pound { "£" }
        .jamaica_dollar { "J$" }
        .jersey_pound { "£" }
        .koruna { "Kč" }
        .kip { "₭" }
        .kuna { "kn" }
        .kyrgyzstan_som { "лв" }
        .lebanon_pound { "£" }
        .lek { "Lek" }
        .lempira { "L" }
        .leu { "lei" }
        .lev { "лв" }
        .liberia_dollar { "\$" }
        .lira { "₺" }
        .azerbaijan_manat { "₼" }
        .mauritius_rupee { "₨" }
        .mexico_peso { "\$" }
        .metical { "MT" }
        .naira { "₦" }
        .namibia_dollar { "\$" }
        .nepal_rupee { "₨" }
        .netherlands_antilles_guilder { "ƒ" }
        .new_taiwan_dollar { "NT$" }
        .new_zealand_dollar { "\$" }
        .north_korea_won { "₩" }
        .norway_krone { "kr" }
        .oman_riyal { "﷼" }
        .pakistan_rupee { "₨" }
        .philipine_peso { "₱" }
        .pula { "P" }
        .qatar_riyal { "﷼" }
        .quetzal { "Q" }
        .rand { "R" }
        .real { "R$" }
        .riel { "៛" }
        .ringgit { "RM" }
        .rupiah { "Rp" }
        .russia_ruble { "₽" }
        .saint_helena_pound { "£" }
        .saudi_arabia_riyal { "﷼" }
        .serbia_dinar { "Дин." }
        .seychelles_rupee { "₨" }
        .shekel { "₪" }
        .shilling { "KSh" }
        .singapore_dollar { "\$" }
        .sol { "S/." }
        .solomon_islands_dollar { "\$" }
        .south_korea_won { "₩" }
        .sri_lanka_rupee { "₨" }
        .suriname_dollar { "\$" }
        .sweden_krona { "kr" }
        .switzerland_franc { "CHF" }
        .syria_pound { "£" }
        .tenge { "₸" }
        .trinidad_and_tobago_dollar { "TT$" }
        .tughrik { "₮" }
        .turkmenistan_manat { "T" }
        .tuvalu_dollar { "\$" }
        .united_kingdom_pound { "£" }
        .united_states_dollar { "\$" }
        .uruguay_peso { "\$U" }
        .uzbekistan_som { "лв" }
        .yen { "¥" }
        .yemen_riyal { "﷼" }
        .yuan { "¥" }
        .zimbabwe_dollar { "Z$" }
        .zloty { "zł" }
    }
}
