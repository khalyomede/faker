module faker

pub struct FakerCountryCodeParameters {
    pub:
        format CountryCodeFormat
}
