module faker

pub struct FakerI64BetweenParameters {
    pub:
        min i64
        max i64
}
