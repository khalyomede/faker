module faker

pub struct FakerF64BetweenParameters {
    pub:
        min f64
        max f64
}
