module faker

pub fn Currency.cases() []Currency {
    return [
        .afghani
        .argentina_peso
        .aruba_guilder
        .australia_dollar
        .azerbaijan_manat
        .bahamas_dollar
        .baht
        .balboa
        .barbados_dollar
        .belarus_ruble
        .belize_dollar
        .bermuda_dollar
        .brunei_darusalam_dollar
        .bolivar
        .boliviano
        .convertible_mark
        .canada_dollar
        .cayman_islands_dollar
        .cedi
        .chile_peso
        .colombia_peso
        .cordoba
        .costa_rica_colon
        .cuba_peso
        .denar
        .denmark_krone
        .dong
        .dominican_republic_peso
        .east_caribbean_dollar
        .egypt_pound
        .euro
        .falkland_islands_pound
        .forint
        .fiji_dollar
        .gibraltar_pound
        .guarani
        .guernsey_pound
        .guyana_dollar
        .hong_kong_dollar
        .hryvnia
        .iceland_krona
        .india_rupee
        .iran_riyal
        .isle_of_man_pound
        .jamaica_dollar
        .jersey_pound
        .koruna
        .kip
        .kuna
        .kyrgyzstan_som
        .lebanon_pound
        .lek
        .lempira
        .leu
        .lev
        .liberia_dollar
        .lira
        .mauritius_rupee
        .mexico_peso
        .metical
        .naira
        .namibia_dollar
        .nepal_rupee
        .netherlands_antilles_guilder
        .new_taiwan_dollar
        .new_zealand_dollar
        .north_korea_won
        .norway_krone
        .oman_riyal
        .pakistan_rupee
        .philipine_peso
        .pula
        .qatar_riyal
        .quetzal
        .rand
        .real
        .riel
        .ringgit
        .rupiah
        .russia_ruble
        .saint_helena_pound
        .saudi_arabia_riyal
        .serbia_dinar
        .seychelles_rupee
        .shekel
        .shilling
        .singapore_dollar
        .sol
        .solomon_islands_dollar
        .south_korea_won
        .sri_lanka_rupee
        .suriname_dollar
        .sweden_krona
        .switzerland_franc
        .syria_pound
        .tenge
        .trinidad_and_tobago_dollar
        .tughrik
        .turkmenistan_manat
        .tuvalu_dollar
        .united_kingdom_pound
        .united_states_dollar
        .uruguay_peso
        .uzbekistan_som
        .yen
        .yemen_riyal
        .yuan
        .zimbabwe_dollar
        .zloty
    ]
}
