module faker

pub fn (country Country) to_alpha_3() string {
    return match country {
        .afghanistan { "AFG" }
        .albania { "ALB" }
        .algeria { "DZA" }
        .andorra { "AND" }
        .angola { "AGO" }
        .antigua_and_barbuda { "ATG" }
        .argentina { "ARG" }
        .armenia { "ARM" }
        .australia { "AUS" }
        .austria { "AUT" }
        .azerbaijan { "AZE" }
        .bahamas { "BHS" }
        .bahrain { "BHR" }
        .bangladesh { "BGD" }
        .barbados { "BRB" }
        .belarus { "BLR" }
        .belgium { "BEL" }
        .belize { "BLZ" }
        .benin { "BEN" }
        .bhutan { "BTN" }
        .bolivia { "BOL" }
        .bosnia_and_herzegovina { "BIH" }
        .botswana { "BWA" }
        .brazil { "BRA" }
        .brunei { "BRN" }
        .bulgaria { "BGR" }
        .burkina_faso { "BFA" }
        .burundi { "BDI" }
        .cabo_verde { "CPV" }
        .cambodia { "KHM" }
        .cameroon { "CMR" }
        .canada { "CAN" }
        .central_african_republic { "CAF" }
        .chad { "TCD" }
        .chile { "CHL" }
        .china { "CHN" }
        .colombia { "COL" }
        .comoros { "COM" }
        .congo { "COG" }
        .costa_rica { "CRI" }
        .croatia { "HRV" }
        .cuba { "CUB" }
        .cyprus { "CYP" }
        .czech_republic { "CZE" }
        .democratic_republic_of_the_congo { "COD" }
        .denmark { "DNK" }
        .djibouti { "DJI" }
        .dominica { "DMA" }
        .dominican_republic { "DOM" }
        .ecuador { "ECU" }
        .egypt { "EGY" }
        .el_salvador { "SLV" }
        .equatorial_guinea { "GNQ" }
        .eritrea { "ERI" }
        .estonia { "EST" }
        .eswatini { "SWZ" }
        .ethiopia { "ETH" }
        .fiji { "FJI" }
        .finland { "FIN" }
        .france { "FRA" }
        .gabon { "GAB" }
        .gambia { "GMB" }
        .georgia { "GEO" }
        .germany { "DEU" }
        .ghana { "GHA" }
        .greece { "GRC" }
        .grenada { "GRD" }
        .guatemala { "GTM" }
        .guinea { "GIN" }
        .guinea_bissau { "GNB" }
        .guyana { "GUY" }
        .haiti { "HTI" }
        .holy_see { "VAT" }
        .honduras { "HND" }
        .hungary { "HUN" }
        .iceland { "ISL" }
        .india { "IND" }
        .indonesia { "IDN" }
        .iran { "IRN" }
        .iraq { "IRQ" }
        .ireland { "IRL" }
        .israel { "ISR" }
        .italy { "ITA" }
        .ivory_coast { "CIV" }
        .jamaica { "JAM" }
        .japan { "JPN" }
        .jordan { "JOR" }
        .kazakhstan { "KAZ" }
        .kenya { "KEN" }
        .kiribati { "KIR" }
        .kosovo { "XKX" }
        .kuwait { "KWT" }
        .kyrgyzstan { "KGZ" }
        .laos { "LAO" }
        .latvia { "LVA" }
        .lebanon { "LBN" }
        .lesotho { "LSO" }
        .liberia { "LBR" }
        .libya { "LBY" }
        .liechtenstein { "LIE" }
        .lithuania { "LTU" }
        .luxembourg { "LUX" }
        .madagascar { "MDG" }
        .malawi { "MWI" }
        .malaysia { "MYS" }
        .maldives { "MDV" }
        .mali { "MLI" }
        .malta { "MLT" }
        .marshall_islands { "MHL" }
        .mauritania { "MRT" }
        .mauritius { "MUS" }
        .mexico { "MEX" }
        .micronesia { "FSM" }
        .moldova { "MDA" }
        .monaco { "MCO" }
        .mongolia { "MNG" }
        .montenegro { "MNE" }
        .morocco { "MAR" }
        .mozambique { "MOZ" }
        .myanmar { "MMR" }
        .namibia { "NAM" }
        .nauru { "NRU" }
        .nepal { "NPL" }
        .netherlands { "NLD" }
        .new_zealand { "NZL" }
        .nicaragua { "NIC" }
        .niger { "NER" }
        .nigeria { "NGA" }
        .north_korea { "PRK" }
        .north_macedonia { "MKD" }
        .norway { "NOR" }
        .oman { "OMN" }
        .pakistan { "PAK" }
        .palau { "PLW" }
        .palestine { "PSE" }
        .panama { "PAN" }
        .papua_new_guinea { "PNG" }
        .paraguay { "PRY" }
        .peru { "PER" }
        .philippines { "PHL" }
        .poland { "POL" }
        .portugal { "PRT" }
        .qatar { "QAT" }
        .romania { "ROU" }
        .russia { "RUS" }
        .rwanda { "RWA" }
        .saint_kitts_and_nevis { "KNA" }
        .saint_lucia { "LCA" }
        .saint_vincent_and_the_grenadines { "VCT" }
        .samoa { "WSM" }
        .san_marino { "SMR" }
        .sao_tome_and_principe { "STP" }
        .saudi_arabia { "SAU" }
        .senegal { "SEN" }
        .serbia { "SRB" }
        .seychelles { "SYC" }
        .sierra_leone { "SLE" }
        .singapore { "SGP" }
        .slovakia { "SVK" }
        .slovenia { "SVN" }
        .solomon_islands { "SLB" }
        .somalia { "SOM" }
        .south_africa { "ZAF" }
        .south_korea { "KOR" }
        .south_sudan { "SSD" }
        .spain { "ESP" }
        .sri_lanka { "LKA" }
        .sudan { "SDN" }
        .suriname { "SUR" }
        .sweden { "SWE" }
        .switzerland { "CHE" }
        .syria { "SYR" }
        .taiwan { "TWN" }
        .tajikistan { "TJK" }
        .tanzania { "TZA" }
        .thailand { "THA" }
        .timor_leste { "TLS" }
        .togo { "TGO" }
        .tonga { "TON" }
        .trinidad_and_tobago { "TTO" }
        .tunisia { "TUN" }
        .turkey { "TUR" }
        .turkmenistan { "TKM" }
        .tuvalu { "TUV" }
        .uganda { "UGA" }
        .ukraine { "UKR" }
        .united_arab_emirates { "ARE" }
        .united_kingdom { "GBR" }
        .united_states { "USA" }
        .uruguay { "URY" }
        .uzbekistan { "UZB" }
        .vanuatu { "VUT" }
        .venezuela { "VEN" }
        .vietnam { "VNM" }
        .yemen { "YEM" }
        .zambia { "ZMB" }
        .zimbabwe { "ZWE" }
    }
}
