module faker

pub struct FakerI16BetweenParameters {
    pub:
        min i16
        max i16
}
