module faker

pub struct FakerI8BetweenParameters {
    pub:
        min i8
        max i8
}
