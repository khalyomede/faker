module faker

pub fn Country.cases() []Country {
    return [
        Country.afghanistan
        Country.albania
        Country.algeria
        Country.andorra
        Country.angola
        Country.antigua_and_barbuda
        Country.argentina
        Country.armenia
        Country.australia
        Country.austria
        Country.azerbaijan
        Country.bahamas
        Country.bahrain
        Country.bangladesh
        Country.barbados
        Country.belarus
        Country.belgium
        Country.belize
        Country.benin
        Country.bhutan
        Country.bolivia
        Country.bosnia_and_herzegovina
        Country.botswana
        Country.brazil
        Country.brunei
        Country.bulgaria
        Country.burkina_faso
        Country.burundi
        Country.cabo_verde
        Country.cambodia
        Country.cameroon
        Country.canada
        Country.central_african_republic
        Country.chad
        Country.chile
        Country.china
        Country.colombia
        Country.comoros
        Country.congo
        Country.costa_rica
        Country.croatia
        Country.cuba
        Country.cyprus
        Country.czech_republic
        Country.democratic_republic_of_the_congo
        Country.denmark
        Country.djibouti
        Country.dominica
        Country.dominican_republic
        Country.ecuador
        Country.egypt
        Country.el_salvador
        Country.equatorial_guinea
        Country.eritrea
        Country.estonia
        Country.eswatini
        Country.ethiopia
        Country.fiji
        Country.finland
        Country.france
        Country.gabon
        Country.gambia
        Country.georgia
        Country.germany
        Country.ghana
        Country.greece
        Country.grenada
        Country.guatemala
        Country.guinea
        Country.guinea_bissau
        Country.guyana
        Country.haiti
        Country.holy_see
        Country.honduras
        Country.hungary
        Country.iceland
        Country.india
        Country.indonesia
        Country.iran
        Country.iraq
        Country.ireland
        Country.israel
        Country.italy
        Country.ivory_coast
        Country.jamaica
        Country.japan
        Country.jordan
        Country.kazakhstan
        Country.kenya
        Country.kiribati
        Country.kosovo
        Country.kuwait
        Country.kyrgyzstan
        Country.laos
        Country.latvia
        Country.lebanon
        Country.lesotho
        Country.liberia
        Country.libya
        Country.liechtenstein
        Country.lithuania
        Country.luxembourg
        Country.madagascar
        Country.malawi
        Country.malaysia
        Country.maldives
        Country.mali
        Country.malta
        Country.marshall_islands
        Country.mauritania
        Country.mauritius
        Country.mexico
        Country.micronesia
        Country.moldova
        Country.monaco
        Country.mongolia
        Country.montenegro
        Country.morocco
        Country.mozambique
        Country.myanmar
        Country.namibia
        Country.nauru
        Country.nepal
        Country.netherlands
        Country.new_zealand
        Country.nicaragua
        Country.niger
        Country.nigeria
        Country.north_korea
        Country.north_macedonia
        Country.norway
        Country.oman
        Country.pakistan
        Country.palau
        Country.palestine
        Country.panama
        Country.papua_new_guinea
        Country.paraguay
        Country.peru
        Country.philippines
        Country.poland
        Country.portugal
        Country.qatar
        Country.romania
        Country.russia
        Country.rwanda
        Country.saint_kitts_and_nevis
        Country.saint_lucia
        Country.saint_vincent_and_the_grenadines
        Country.samoa
        Country.san_marino
        Country.sao_tome_and_principe
        Country.saudi_arabia
        Country.senegal
        Country.serbia
        Country.seychelles
        Country.sierra_leone
        Country.singapore
        Country.slovakia
        Country.slovenia
        Country.solomon_islands
        Country.somalia
        Country.south_africa
        Country.south_korea
        Country.south_sudan
        Country.spain
        Country.sri_lanka
        Country.sudan
        Country.suriname
        Country.sweden
        Country.switzerland
        Country.syria
        Country.taiwan
        Country.tajikistan
        Country.tanzania
        Country.thailand
        Country.timor_leste
        Country.togo
        Country.tonga
        Country.trinidad_and_tobago
        Country.tunisia
        Country.turkey
        Country.turkmenistan
        Country.tuvalu
        Country.uganda
        Country.ukraine
        Country.united_arab_emirates
        Country.united_kingdom
        Country.united_states
        Country.uruguay
        Country.uzbekistan
        Country.vanuatu
        Country.venezuela
        Country.vietnam
        Country.yemen
        Country.zambia
        Country.zimbabwe
    ]
}
