module faker

pub enum CountryCodeFormat {
    alpha_2
    alpha_3
}
