module faker

pub struct FakerU32BetweenParameters {
    pub:
        min u32
        max u32
}
