module faker

pub fn (country Country) to_alpha_2() string {
    return match country {
        .afghanistan { "AF" }
        .albania { "AL" }
        .algeria { "DZ" }
        .andorra { "AD" }
        .angola { "AO" }
        .antigua_and_barbuda { "AG" }
        .argentina { "AR" }
        .armenia { "AM" }
        .australia { "AU" }
        .austria { "AT" }
        .azerbaijan { "AZ" }
        .bahamas { "BS" }
        .bahrain { "BH" }
        .bangladesh { "BD" }
        .barbados { "BB" }
        .belarus { "BY" }
        .belgium { "BE" }
        .belize { "BZ" }
        .benin { "BJ" }
        .bhutan { "BT" }
        .bolivia { "BO" }
        .bosnia_and_herzegovina { "BA" }
        .botswana { "BW" }
        .brazil { "BR" }
        .brunei { "BN" }
        .bulgaria { "BG" }
        .burkina_faso { "BF" }
        .burundi { "BI" }
        .cabo_verde { "CV" }
        .cambodia { "KH" }
        .cameroon { "CM" }
        .canada { "CA" }
        .central_african_republic { "CF" }
        .chad { "TD" }
        .chile { "CL" }
        .china { "CN" }
        .colombia { "CO" }
        .comoros { "KM" }
        .congo { "CG" }
        .costa_rica { "CR" }
        .croatia { "HR" }
        .cuba { "CU" }
        .cyprus { "CY" }
        .czech_republic { "CZ" }
        .democratic_republic_of_the_congo { "CD" }
        .denmark { "DK" }
        .djibouti { "DJ" }
        .dominica { "DM" }
        .dominican_republic { "DO" }
        .ecuador { "EC" }
        .egypt { "EG" }
        .el_salvador { "SV" }
        .equatorial_guinea { "GQ" }
        .eritrea { "ER" }
        .estonia { "EE" }
        .eswatini { "SZ" }
        .ethiopia { "ET" }
        .fiji { "FJ" }
        .finland { "FI" }
        .france { "FR" }
        .gabon { "GA" }
        .gambia { "GM" }
        .georgia { "GE" }
        .germany { "DE" }
        .ghana { "GH" }
        .greece { "GR" }
        .grenada { "GD" }
        .guatemala { "GT" }
        .guinea { "GN" }
        .guinea_bissau { "GW" }
        .guyana { "GY" }
        .haiti { "HT" }
        .holy_see { "VA" }
        .honduras { "HN" }
        .hungary { "HU" }
        .iceland { "IS" }
        .india { "IN" }
        .indonesia { "ID" }
        .iran { "IR" }
        .iraq { "IQ" }
        .ireland { "IE" }
        .israel { "IL" }
        .italy { "IT" }
        .ivory_coast { "CI" }
        .jamaica { "JM" }
        .japan { "JP" }
        .jordan { "JO" }
        .kazakhstan { "KZ" }
        .kenya { "KE" }
        .kiribati { "KI" }
        .kosovo { "XK" }
        .kuwait { "KW" }
        .kyrgyzstan { "KG" }
        .laos { "LA" }
        .latvia { "LV" }
        .lebanon { "LB" }
        .lesotho { "LS" }
        .liberia { "LR" }
        .libya { "LY" }
        .liechtenstein { "LI" }
        .lithuania { "LT" }
        .luxembourg { "LU" }
        .madagascar { "MG" }
        .malawi { "MW" }
        .malaysia { "MY" }
        .maldives { "MV" }
        .mali { "ML" }
        .malta { "MT" }
        .marshall_islands { "MH" }
        .mauritania { "MR" }
        .mauritius { "MU" }
        .mexico { "MX" }
        .micronesia { "FM" }
        .moldova { "MD" }
        .monaco { "MC" }
        .mongolia { "MN" }
        .montenegro { "ME" }
        .morocco { "MA" }
        .mozambique { "MZ" }
        .myanmar { "MM" }
        .namibia { "NA" }
        .nauru { "NR" }
        .nepal { "NP" }
        .netherlands { "NL" }
        .new_zealand { "NZ" }
        .nicaragua { "NI" }
        .niger { "NE" }
        .nigeria { "NG" }
        .north_korea { "KP" }
        .north_macedonia { "MK" }
        .norway { "NO" }
        .oman { "OM" }
        .pakistan { "PK" }
        .palau { "PW" }
        .palestine { "PS" }
        .panama { "PA" }
        .papua_new_guinea { "PG" }
        .paraguay { "PY" }
        .peru { "PE" }
        .philippines { "PH" }
        .poland { "PL" }
        .portugal { "PT" }
        .qatar { "QA" }
        .romania { "RO" }
        .russia { "RU" }
        .rwanda { "RW" }
        .saint_kitts_and_nevis { "KN" }
        .saint_lucia { "LC" }
        .saint_vincent_and_the_grenadines { "VC" }
        .samoa { "WS" }
        .san_marino { "SM" }
        .sao_tome_and_principe { "ST" }
        .saudi_arabia { "SA" }
        .senegal { "SN" }
        .serbia { "RS" }
        .seychelles { "SC" }
        .sierra_leone { "SL" }
        .singapore { "SG" }
        .slovakia { "SK" }
        .slovenia { "SI" }
        .solomon_islands { "SB" }
        .somalia { "SO" }
        .south_africa { "ZA" }
        .south_korea { "KR" }
        .south_sudan { "SS" }
        .spain { "ES" }
        .sri_lanka { "LK" }
        .sudan { "SD" }
        .suriname { "SR" }
        .sweden { "SE" }
        .switzerland { "CH" }
        .syria { "SY" }
        .taiwan { "TW" }
        .tajikistan { "TJ" }
        .tanzania { "TZ" }
        .thailand { "TH" }
        .timor_leste { "TL" }
        .togo { "TG" }
        .tonga { "TO" }
        .trinidad_and_tobago { "TT" }
        .tunisia { "TN" }
        .turkey { "TR" }
        .turkmenistan { "TM" }
        .tuvalu { "TV" }
        .uganda { "UG" }
        .ukraine { "UA" }
        .united_arab_emirates { "AE" }
        .united_kingdom { "GB" }
        .united_states { "US" }
        .uruguay { "UY" }
        .uzbekistan { "UZ" }
        .vanuatu { "VU" }
        .venezuela { "VE" }
        .vietnam { "VN" }
        .yemen { "YE" }
        .zambia { "ZM" }
        .zimbabwe { "ZW" }
    }
}
