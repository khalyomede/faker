module faker

pub struct FakerU16BetweenParameters {
    pub:
        min u16
        max u16
}
